module top_tb;

fifo_tb dut();
scfifo_tb dut2();
endmodule